// top level testbench
// in order to run must set the input matrix
// then reset and let the input be read in one pixel at a time
// to run it again would just need to adjust what the input matrix is
// you do not need to reset it   
          
module convNN_top_test(); 
	parameter filtDimension = 3, bitWidth =4, inputWidth = 8, weightWidth = 18, biasWidth = 2, outputSize = 10, 
	numFilt = 2;
	
	logic clk_p, clk_n, reset;
	logic signed [bitWidth-1:0] inputPixel;
	logic signed [bitWidth-1:0] copyOutputDL [outputSize-1:0];
	logic signed [bitWidth-1:0] outputSoftmax [outputSize-1:0];
	
	logic signed [bitWidth-1:0] inputMatrix [63:0];
	logic outputValid;
	
//    assign inputMatrix = {
//    16'd0, 16'd0, 16'd0, 16'd0, 16'd0, 16'd0, 16'd0, 16'd0,
//    16'd1, 16'd1, 16'd1, 16'd1, 16'd1, 16'd1, 16'd1 ,16'd1,
//    16'd2, 16'd2, 16'd2, 16'd2, 16'd2, 16'd2, 16'd2, 16'd2,
//    16'd3, 16'd3, 16'd3, 16'd3, 16'd3, 16'd3, 16'd3 ,16'd3,
//    16'd4, 16'd4, 16'd4, 16'd4, 16'd4, 16'd4, 16'd4 ,16'd4,
//    16'd5, 16'd5, 16'd5, 16'd5, 16'd5, 16'd5, 16'd5, 16'd5,
//    16'd6, 16'd6, 16'd6, 16'd6, 16'd6, 16'd6, 16'd6 ,16'd6,
//    16'd7, 16'd7, 16'd7, 16'd7, 16'd7, 16'd7, 16'd7 ,16'd7
//    };
    
//    assign inputMatrix = {
//    17'b00001000000000000, 17'd0, 17'd0, 17'd0, 17'd0, 17'd0, 17'd0, 17'd0,
//    17'd0, 17'b00001000000000000, 17'd0, 17'd0, 17'd0, 17'd0, 17'd0, 17'd0,
//    17'd0, 17'd0, 17'b00001000000000000, 17'd0, 17'd0, 17'd0, 17'd0, 17'd0,
//    17'd0, 17'd0, 17'd0, 17'b00001000000000000, 17'd0, 17'd0, 17'd0, 17'd0,
//    17'd0, 17'd0, 17'd0, 17'd0, 17'b00001000000000000, 17'd0, 17'd0, 17'd0,
//    17'd0, 17'd0, 17'd0, 17'd0, 17'd0, 17'b00001000000000000, 17'd0, 17'd0,
//    17'd0, 17'd0, 17'd0, 17'd0, 17'd0, 17'd0, 17'b00001000000000000, 17'd0,
//    17'd0, 17'd0, 17'd0, 17'd0, 17'd0, 17'd0, 17'd0, 17'b00001000000000000
//    };
	
//	assign inputMatrix = {
//    17'b00001000000000000, 17'b00001000000000000, 17'b00001000000000000, 17'b00001000000000000, 17'b00001000000000000,17'b00001000000000000, 17'b00001000000000000, 17'b00001000000000000,
//    17'b00001000000000000, 17'b00001000000000000, 17'b00001000000000000, 17'b00001000000000000, 17'b00001000000000000,17'b00001000000000000, 17'b00001000000000000, 17'b00001000000000000,
//    17'b00001000000000000, 17'b00001000000000000, 17'b00001000000000000, 17'b00001000000000000, 17'b00001000000000000,17'b00001000000000000, 17'b00001000000000000, 17'b00001000000000000,
//    17'b00001000000000000, 17'b00001000000000000, 17'b00001000000000000, 17'b00001000000000000, 17'b00001000000000000,17'b00001000000000000, 17'b00001000000000000, 17'b00001000000000000,
//    17'b00001000000000000, 17'b00001000000000000, 17'b00001000000000000, 17'b00001000000000000, 17'b00001000000000000,17'b00001000000000000, 17'b00001000000000000, 17'b00001000000000000,
//    17'b00001000000000000, 17'b00001000000000000, 17'b00001000000000000, 17'b00001000000000000, 17'b00001000000000000,17'b00001000000000000, 17'b00001000000000000, 17'b00001000000000000,
//    17'b00001000000000000, 17'b00001000000000000, 17'b00001000000000000, 17'b00001000000000000, 17'b00001000000000000,17'b00001000000000000, 17'b00001000000000000, 17'b00001000000000000,
//    17'b00001000000000000, 17'b00001000000000000, 17'b00001000000000000, 17'b00001000000000000, 17'b00001000000000000,17'b00001000000000000, 17'b00001000000000000, 17'b00001000000000000
//    };


//assign inputMatrix = {
//    16'b0000000010011100, 16'b0000000110001111, 16'b0000000001111101, 16'b1111111110110011, 16'b1111111101111101, 16'b0000000001000101, 16'b0000000010011100, 16'b0000000011001010,
//    16'b1111111010010110, 16'b0000000010111101, 16'b0000000111100000, 16'b1111111111111001, 16'b0000000100101001, 16'b1111111110101111, 16'b0000000000111011, 16'b0000000000100010,
//    16'b0000000010011100, 16'b0000000110001111, 16'b0000000001111101, 16'b1111111110110011, 16'b1111111101111101, 16'b0000000001000101, 16'b0000000010011100, 16'b0000000011001010,
//    16'b1111111010010110, 16'b0000000010111101, 16'b0000000111100000, 16'b1111111111111001, 16'b0000000100101001, 16'b1111111110101111, 16'b0000000000111011, 16'b0000000000100010,
//    16'b0000000010011100, 16'b0000000110001111, 16'b0000000001111101, 16'b1111111110110011, 16'b1111111101111101, 16'b0000000001000101, 16'b0000000010011100, 16'b0000000011001010,
//    16'b1111111010010110, 16'b0000000010111101, 16'b0000000111100000, 16'b1111111111111001, 16'b0000000100101001, 16'b1111111110101111, 16'b0000000000111011, 16'b0000000000100010,
//    16'b0000000010011100, 16'b0000000110001111, 16'b0000000001111101, 16'b1111111110110011, 16'b1111111101111101, 16'b0000000001000101, 16'b0000000010011100, 16'b0000000011001010,
//    16'b1111111010010110, 16'b0000000010111101, 16'b0000000111100000, 16'b1111111111111001, 16'b0000000100101001, 16'b1111111110101111, 16'b0000000000111011, 16'b0000000000100010
//    };
    assign inputMatrix = {
    17'd0, 17'd0, 17'd0, 17'd0, 17'd0, 17'd0, 17'd0, 17'd0,
    17'd1, 17'd1, 17'd1, 17'd1, 17'd1, 17'd1, 17'd1, 17'd1,
    17'd2, 17'd2, 17'd2, 17'd2, 17'd2, 17'd2, 17'd2, 17'd2,
    17'd3, 17'd3, 17'd3, 17'd3, 17'd3, 17'd3, 17'd3, 17'd3,
    17'd4, 17'd4, 17'd4, 17'd4, 17'd4, 17'd4, 17'd4, 17'd4,
    17'd5, 17'd5, 17'd5, 17'd5, 17'd5, 17'd5, 17'd5, 17'd5,
    17'd6, 17'd6, 17'd6, 17'd6, 17'd6, 17'd6, 17'd6, 17'd6,
    17'd7, 17'd7, 17'd7, 17'd7, 17'd7, 17'd7, 17'd7, 17'd7
    };
	conv2d_connector #(3,4,8,18,2,10,2,2) dut (.*);
	
	// Set up a simulated clock.
	parameter CLOCK_PERIOD=100;
	initial begin
        clk_p <= 0;
        clk_n <= 1;
        forever #(CLOCK_PERIOD/2) begin
            clk_p <= ~clk_p;
            clk_n <= ~clk_n;
        end
    end
	integer i,j;
	
	
	
	initial begin
	reset <= 1; 
	//inputPixel <= 16'b0001000000000000;@(posedge clk_p);
	
	 //inputPixel <= inputMatrix[63]; @(posedge clk_p);
	 inputPixel <= 10'd2; @(posedge clk_p);
	 
	 for(int i =62; i>=0; i--) begin
	  // reset <= 0; inputPixel <= inputMatrix[i]; @(posedge clk_p);
	  reset<=0; inputPixel <= 10'd2; @(posedge clk_p);
	 end

	 repeat(300) @(posedge clk_p);

	 // inputPixel <= 18'd6; repeat(100) @(posedge clk_p);
	   
	  //inputPixel <= 17'b00001000000000000; repeat(64)@(posedge clk_p);
	  
	  for(i=0; i<128; i++)begin
	  $display("%b", dut.dense.denseSums[0].sumColumns.sums.input_data[i]);
	   end @(posedge clk_p);
	
	$stop; // End the simulation.
	end
endmodule
	